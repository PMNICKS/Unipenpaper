�PNG

   IHDR   �   �   ��6   �PLTE����((   �::�%%�����������������  ���������222����  �00���,,,===������������EEE�����������iiiii!!!rrr�NNN����������bb�}}����\\��������uu�EE�MM^^^)�я  �IDATx��	S�8F�J��dْ����̂��ۖaj�YrM-���WE��"j_� � � � bf��yj������S;������д׫�js�pj��X��h���ʈ�F��:��"E������(Zm�����@~Jc��N�so�}�� ��?�1ګ��S;���hy��9;��>~����t{j�=�[ڗ�ż��{�X�V�s�������|�[�}��ק���Vi��fd�4F��f�G����F{�4f��i~W��gyҺ_�}=���}8w���}9<�gϋ�f�<@�G��������s��Kk_�T�������|;$��.������̤Q{y��j�N/~/������#�ў�4��>��������~�7Wi�z�-#�Ɠ�����G��)�#��b����a<��OM��r+�� o!|�ܬ�:�f�'�-��o�xS=��>(
�\�?|����N8H%��@!�
p��O@��� Ȇ89�A�A��� � � � � � �$,@H�� ��b��6cZ�R+d�
Y1W��sݲF�8G"�eѕ�5R���g�]^r.j�%w�q.��\�,�u�L�����ꎕB$,w~C�͙��H��`�aDlF�)Q�X�eL�4Nuu�5$.�PYi��N�r�q��tp���@I92�+�9ܜL��dJnZ���2�R�P@�
�s�0�M���ƈ�d#��/3hm�ƾe=4�)�t�4mc�5E����TI<�]�%PY���i�\�V�R�y�jlWax.����k�uJ�ܽ�/�2���2R�JGK�u�+��
_T�*�[��֠̋4~�b�*��Jk��6Z��(�10�����(\(�q��t����N��z�jИ@kƪ��s�F��-++�����Y	�t-���L�c�i��F4�Su'=��i\�H�8jPqik���[��M�
3X�%�^�Ôi�GҖ� ���T^�fZb~Jc�h��5Nq�~�!�M-�g��{�un�({Y��$��J�'=+]e}�g?:Ӆ�u���c���çJ��l+�KY!�/-�b|j���("�t�Racm�o;�um6}�M{,{�����YW��Gi��X�����G��[J�nZ�Lk�0��$�U��o���,��%4H��R�o��� �    IEND�B`�