�PNG

   IHDR   �   �   ���   lPLTE���    �����������Ǘ��  ���+,+%'%787���	���]^]121MMM��ស�BCB���=>=llk���������VVUѶ�  �IDATx��mo�0��!�N���������4�����p�gO~�G�3�B��@ ���.�w�5<c����[g��T�T�JP�V�p�o)�ԺT_�ɷ�5�f��޷�eg�����,�i�-R9�Yf͏I�>��#"m�[����-b^2���|+Z ����$]�[��"v�q�s-"۝k�8)��y&�B�d�av#N���"��9YB�Mk�����b�8I!�H')�E��"�Hf��}+Z k�ݐ�X�Z����Z�� �Z�$��k�n��x��[D-*��_�5KKs�r )�ݐ��)�բA����j%��"jQ­��ZH�C-�#xN��oEd��;�Z4�Hz
R�%�a;~��iN^i70�v�r�$���i�����cg�Dba�1*�oO�E�����R����|�;h�S�.๼D[�>Ls�&f\���[M�>p�S�ğ�Y�7T���0�EΧi���U������x`p$���ŷ�EMdV=���y�4=f��1���17�Bs�:a��&�+	�de)f��2���eIM�����&3݁��˲C�rc:+K��'$L��B�eY�0����<7����RJnb�do����t1e�J0��dt��)�,A�9TBVHDn�lPs�l�=`N����w'$�M�	��BM�w!'$V����f	��f�WȽ�ֳY��rZ���o5��0]�Ŭ3�d�y��Ilo���r��!Y��IE�C3cV9�݁@ ��*�I_4��ch    IEND�B`�